///////////////////////////////////////////////////////////////////////////////
// BEGIN Global Parameters
///////////////////////////////////////////////////////////////////////////////
localparam G_AXI_AWADDR_INDEX   = 0;
localparam G_AXI_AWADDR_WIDTH   = C_AXI_ADDR_WIDTH;
localparam G_AXI_AWPROT_INDEX   = G_AXI_AWADDR_INDEX + G_AXI_AWADDR_WIDTH;
localparam G_AXI_AWPROT_WIDTH   = 3;
localparam G_AXI_AWSIZE_INDEX   = G_AXI_AWPROT_INDEX + G_AXI_AWPROT_WIDTH;
localparam G_AXI_AWSIZE_WIDTH   = (C_AXI_PROTOCOL == 2) ? 0 : 3;
localparam G_AXI_AWBURST_INDEX  = G_AXI_AWSIZE_INDEX + G_AXI_AWSIZE_WIDTH;
localparam G_AXI_AWBURST_WIDTH  = (C_AXI_PROTOCOL == 2) ? 0 : 2;
localparam G_AXI_AWCACHE_INDEX  = G_AXI_AWBURST_INDEX + G_AXI_AWBURST_WIDTH;
localparam G_AXI_AWCACHE_WIDTH  = (C_AXI_PROTOCOL == 2) ? 0 : 4;
localparam G_AXI_AWLEN_INDEX    = G_AXI_AWCACHE_INDEX + G_AXI_AWCACHE_WIDTH;
localparam G_AXI_AWLEN_WIDTH    = (C_AXI_PROTOCOL == 2) ? 0 : (C_AXI_PROTOCOL == 1) ? 4 : 8;
localparam G_AXI_AWLOCK_INDEX   = G_AXI_AWLEN_INDEX + G_AXI_AWLEN_WIDTH;
localparam G_AXI_AWLOCK_WIDTH   = (C_AXI_PROTOCOL == 2) ? 0 : (C_AXI_PROTOCOL == 1) ? 2 : 1;
localparam G_AXI_AWID_INDEX     = G_AXI_AWLOCK_INDEX + G_AXI_AWLOCK_WIDTH;
localparam G_AXI_AWID_WIDTH     = (C_AXI_PROTOCOL == 2) ? 0 : C_AXI_ID_WIDTH;
localparam G_AXI_AWQOS_INDEX    = G_AXI_AWID_INDEX + G_AXI_AWID_WIDTH;
localparam G_AXI_AWQOS_WIDTH    = (C_AXI_PROTOCOL == 2) ? 0 : 4;
localparam G_AXI_AWREGION_INDEX = G_AXI_AWQOS_INDEX + G_AXI_AWQOS_WIDTH;
localparam G_AXI_AWREGION_WIDTH = (C_AXI_PROTOCOL == 2) ? 0 : (C_AXI_SUPPORTS_REGION_SIGNALS == 0) ? 0 : 4;
localparam G_AXI_AWUSER_INDEX   = G_AXI_AWREGION_INDEX + G_AXI_AWREGION_WIDTH;
localparam G_AXI_AWUSER_WIDTH   = (C_AXI_PROTOCOL == 2) ? 0 : (C_AXI_SUPPORTS_USER_SIGNALS == 0) ? 0 : C_AXI_AWUSER_WIDTH;
localparam G_AXI_AWPAYLOAD_WIDTH = G_AXI_AWUSER_INDEX + G_AXI_AWUSER_WIDTH;
localparam G_AXI_ARADDR_INDEX   = 0;
localparam G_AXI_ARADDR_WIDTH   = C_AXI_ADDR_WIDTH;
localparam G_AXI_ARPROT_INDEX   = G_AXI_ARADDR_INDEX + G_AXI_ARADDR_WIDTH;
localparam G_AXI_ARPROT_WIDTH   = 3;
localparam G_AXI_ARSIZE_INDEX   = G_AXI_ARPROT_INDEX + G_AXI_ARPROT_WIDTH;
localparam G_AXI_ARSIZE_WIDTH   = (C_AXI_PROTOCOL == 2) ? 0 : 3;
localparam G_AXI_ARBURST_INDEX  = G_AXI_ARSIZE_INDEX + G_AXI_ARSIZE_WIDTH;
localparam G_AXI_ARBURST_WIDTH  = (C_AXI_PROTOCOL == 2) ? 0 : 2;
localparam G_AXI_ARCACHE_INDEX  = G_AXI_ARBURST_INDEX + G_AXI_ARBURST_WIDTH;
localparam G_AXI_ARCACHE_WIDTH  = (C_AXI_PROTOCOL == 2) ? 0 : 4;
localparam G_AXI_ARLEN_INDEX    = G_AXI_ARCACHE_INDEX + G_AXI_ARCACHE_WIDTH;
localparam G_AXI_ARLEN_WIDTH    = (C_AXI_PROTOCOL == 2) ? 0 : (C_AXI_PROTOCOL == 1) ? 4 : 8;
localparam G_AXI_ARLOCK_INDEX   = G_AXI_ARLEN_INDEX + G_AXI_ARLEN_WIDTH;
localparam G_AXI_ARLOCK_WIDTH   = (C_AXI_PROTOCOL == 2) ? 0 : (C_AXI_PROTOCOL == 1) ? 2 : 1;
localparam G_AXI_ARID_INDEX     = G_AXI_ARLOCK_INDEX + G_AXI_ARLOCK_WIDTH;
localparam G_AXI_ARID_WIDTH     = (C_AXI_PROTOCOL == 2) ? 0 : C_AXI_ID_WIDTH;
localparam G_AXI_ARQOS_INDEX    = G_AXI_ARID_INDEX + G_AXI_ARID_WIDTH;
localparam G_AXI_ARQOS_WIDTH    = (C_AXI_PROTOCOL == 2) ? 0 : 4;
localparam G_AXI_ARREGION_INDEX = G_AXI_ARQOS_INDEX + G_AXI_ARQOS_WIDTH;
localparam G_AXI_ARREGION_WIDTH = (C_AXI_PROTOCOL == 2) ? 0 : (C_AXI_SUPPORTS_REGION_SIGNALS == 0) ? 0 : 4;
localparam G_AXI_ARUSER_INDEX   = G_AXI_ARREGION_INDEX + G_AXI_ARREGION_WIDTH;
localparam G_AXI_ARUSER_WIDTH   = (C_AXI_PROTOCOL == 2) ? 0 : (C_AXI_SUPPORTS_USER_SIGNALS == 0) ? 0 : C_AXI_ARUSER_WIDTH;
localparam G_AXI_ARPAYLOAD_WIDTH = G_AXI_ARUSER_INDEX + G_AXI_ARUSER_WIDTH;
// Write channel widths
localparam G_AXI_WDATA_INDEX    = 0;
localparam G_AXI_WDATA_WIDTH    = C_AXI_DATA_WIDTH;
localparam G_AXI_WSTRB_INDEX    = G_AXI_WDATA_INDEX + G_AXI_WDATA_WIDTH;
localparam G_AXI_WSTRB_WIDTH    = C_AXI_DATA_WIDTH / 8;
localparam G_AXI_WLAST_INDEX    = G_AXI_WSTRB_INDEX + G_AXI_WSTRB_WIDTH;
localparam G_AXI_WLAST_WIDTH    = (C_AXI_PROTOCOL == 2) ? 0 : 1;
localparam G_AXI_WID_INDEX      = G_AXI_WLAST_INDEX + G_AXI_WLAST_WIDTH;
localparam G_AXI_WID_WIDTH      = (C_AXI_PROTOCOL != 1) ? 0 : C_AXI_ID_WIDTH;
localparam G_AXI_WUSER_INDEX    = G_AXI_WID_INDEX + G_AXI_WID_WIDTH;
localparam G_AXI_WUSER_WIDTH    = (C_AXI_PROTOCOL == 2) ? 0 : (C_AXI_SUPPORTS_USER_SIGNALS == 0) ? 0 : C_AXI_WUSER_WIDTH;
localparam G_AXI_WPAYLOAD_WIDTH = G_AXI_WUSER_INDEX + G_AXI_WUSER_WIDTH;
// Write Response channel Widths
localparam G_AXI_BRESP_INDEX    = 0;
localparam G_AXI_BRESP_WIDTH    = 2;
localparam G_AXI_BID_INDEX      = G_AXI_BRESP_INDEX + G_AXI_BRESP_WIDTH;
localparam G_AXI_BID_WIDTH      = (C_AXI_PROTOCOL == 2) ? 0 : C_AXI_ID_WIDTH;
localparam G_AXI_BUSER_INDEX    = G_AXI_BID_INDEX + G_AXI_BID_WIDTH;
localparam G_AXI_BUSER_WIDTH    = (C_AXI_PROTOCOL == 2) ? 0 : (C_AXI_SUPPORTS_USER_SIGNALS == 0) ? 0 : C_AXI_BUSER_WIDTH;
localparam G_AXI_BPAYLOAD_WIDTH = G_AXI_BUSER_INDEX + G_AXI_BUSER_WIDTH;
// Read channel widths
localparam G_AXI_RDATA_INDEX    = 0;
localparam G_AXI_RDATA_WIDTH    = C_AXI_DATA_WIDTH;
localparam G_AXI_RRESP_INDEX    = G_AXI_RDATA_INDEX + G_AXI_RDATA_WIDTH;
localparam G_AXI_RRESP_WIDTH    = 2;
localparam G_AXI_RLAST_INDEX    = G_AXI_RRESP_INDEX + G_AXI_RRESP_WIDTH;
localparam G_AXI_RLAST_WIDTH    = (C_AXI_PROTOCOL == 2) ? 0 : 1;
localparam G_AXI_RID_INDEX      = G_AXI_RLAST_INDEX + G_AXI_RLAST_WIDTH;
localparam G_AXI_RID_WIDTH      = (C_AXI_PROTOCOL == 2) ? 0 : C_AXI_ID_WIDTH;
localparam G_AXI_RUSER_INDEX    = G_AXI_RID_INDEX + G_AXI_RID_WIDTH;
localparam G_AXI_RUSER_WIDTH    = (C_AXI_PROTOCOL == 2) ? 0 : (C_AXI_SUPPORTS_USER_SIGNALS == 0) ? 0 : C_AXI_RUSER_WIDTH;
localparam G_AXI_RPAYLOAD_WIDTH = G_AXI_RUSER_INDEX + G_AXI_RUSER_WIDTH;
